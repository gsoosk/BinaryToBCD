library verilog;
use verilog.vl_types.all;
entity binary_into_bcd_with_controller_TB is
end binary_into_bcd_with_controller_TB;
