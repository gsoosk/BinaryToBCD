library verilog;
use verilog.vl_types.all;
entity comb_TB is
end comb_TB;
