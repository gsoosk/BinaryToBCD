library verilog;
use verilog.vl_types.all;
entity counter_TB is
end counter_TB;
